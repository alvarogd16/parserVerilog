module adder #(parameter F = 2, parameter Y=5, H=6)(output x); // #(parameter F = 2, parameter Y=5)(in_a, in_b, out) (input a, in_b, output reg out)

// localparam [N*2:1] A = N;
// localparam hola = "hola";
// localparam number = 5.5;
// localparam number1 = 2'b01;
// localparam number2 = 8'hA5;

// parameter hola = "hola";
// parameter number = 5.5;
// parameter number1 = 2'b01;
// parameter number2 = 8'hA5;

// parameter N = 8, C = 6, G = 4;
// parameter julita = 1;
// parameter [N*2/4-2*(1+1+1):1] B = 8-N, J = 6;

// input in_a, in_b;
// input wire in_c, in_d;
input [16:5] in_e;

// output reg o_a, o_b;
// output wire o_c, o_d;
// output o_e;

// assign out = in_a + in_b;

initial begin
    // $display("N %d %b", N, N);
end

endmodule